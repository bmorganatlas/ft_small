["Quas in recusandae qui explicabo eligendi. Facilis reprehenderit molestiae ut. Porro illo et impedit dolore eos.", "Hic quas ut odit autem dolores voluptatem doloribus. Velit voluptas ipsum. Aspernatur id non numquam ut temporibus sit ut.", "Commodi debitis sit saepe molestias voluptatem. Quis praesentium adipisci iure. Saepe ipsam et provident sit tenetur. Nihil rem sequi saepe ut perferendis pariatur magni. Est dolor odit laboriosam quae aut aperiam consequatur.", "Saepe architecto a qui exercitationem mollitia repudiandae iusto. In corrupti inventore praesentium similique deleniti quidem. Autem quos sint at consectetur distinctio est ex. Alias sed eveniet qui et quam.", "Placeat velit asperiores nostrum qui officia doloribus. Optio sint corporis adipisci. Fugit saepe tempora.", "Soluta impedit enim quam consequatur mollitia. Asperiores autem quas. Quia modi accusamus error deserunt. Veritatis et totam aliquid molestiae sequi distinctio neque."]