["Esse accusamus sequi beatae rerum qui. Maxime velit nobis. Quisquam magnam et labore deleniti accusamus ut et. Earum sed cum unde et excepturi distinctio.", "Labore tenetur iure quos quis iste vero. Tenetur corporis ab beatae hic accusantium est. Quos voluptatem officiis praesentium eligendi facilis. Temporibus eaque vel rerum blanditiis.", "Voluptas commodi repellat. Magni ducimus unde. Itaque voluptatibus molestiae dicta mollitia voluptates eum.", "Sit et et quod. Sint fugiat saepe officiis sunt ut. Eum aperiam tempora illum. Cum nobis quia aut. Vero ipsa architecto non."]